`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:     A*STAR IHPC
// Engineer:    Gerlinghoff Daniel
// Create Date: 18/05/2021
//
// Description: Automatically generated package with config for linear layers
//
//////////////////////////////////////////////////////////////////////////////////


package pkg_linear;
	localparam int LINUNITS = 1;
	localparam int LIN_SIZE = 84;
	localparam int LIN_CHANNELS_MAX = 120;
	localparam int ACT_BITS = 3;
	localparam int WGT_BITS = 3;
	localparam int SUM_BITS = 10;

endpackage
